`timescale 1ns / 1ps

module TOP_VGA #(
  parameter DATA_WIDTH = 16,
  parameter ADDR_WIDTH = 19
 )(
    input  wire        clk,
    input  wire        clk_en,
    input  wire        rst,
    
    // Block RAM Port B (read-only)
    input  wire [7:0]  din,     // BRAM doutb
    output wire        WES,     // Port A write enable
    output wire [7:0]  dout,    // Port A write data
    output wire [18:0] addr,    // BRAM address

    // VGA interface
    output wire [7:0]  rgb,
    output wire        hsyncb,
    output wire        vsyncb,

    // Slide switches
    input  wire [3:0]  sw       // SW[0] : show / hide, SW[3:1] : Y offset
 );

    // ───────────────────────────────
    // Display config / control
    // ───────────────────────────────
    wire [9:0] offset_x;
    wire [8:0] offset_y;
    wire       blank_region;

    wire       img_enable;      // SW[0] = 1 -> show image
    wire [2:0] step_sel;        // SW[3:1] -> Yoffset step

    assign img_enable = sw[0];
    assign step_sel   = sw[3:1];

    localparam XRES = 320;
    localparam YRES = 240;

    // Xoffset = 0, Yoffset = SW[3:1] * 32 pixel
    assign offset_x = 10'd0;
    assign offset_y = {step_sel, 5'b00000};  // step_sel << 5 = *32

    // ───────────────────────────────
    // BRAM -> VGA data path
    // ───────────────────────────────
    wire [7:0]  pixel_raw;       // raw data from BRAM
    wire [7:0]  pixel_masked;    // masked data based on SW[0]
    wire [18:0] mem_rd_addr;     // address generated by VGA

    assign pixel_raw    = din;
    assign pixel_masked = img_enable ? pixel_raw : 8'h00;  // black if SW[0]=0

    // BRAM Port A outputs (unused, constant)
    assign addr = mem_rd_addr;
    assign WES  = 1'b0;
    assign dout = 8'd0;

    // ───────────────────────────────
    // VGA timing + pixel generator
    // ───────────────────────────────
    VGA_module vga (
        .clk        (clk),
        .clk_en     (clk_en),
        .rst        (rst),
        .data       (pixel_masked),
        .hsyncb     (hsyncb),
        .vsyncb     (vsyncb),
        .Xoffset    (offset_x),
        .Yoffset    (offset_y),
        .imageWidth (XRES),
        .imageHeight(YRES),
        .addr       (mem_rd_addr),
        .video_off  (blank_region),
        .rgb        (rgb)
    );

endmodule