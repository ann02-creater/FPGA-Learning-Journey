`timescale 1ns / 1ps

module tb_block_vga();


endmodule
